100 10 0 0 0 0 0 0 0 0 0 0 0 0 0 Jungle 82 0 ph 0 0 1 0 0 100 0